module addressdecoder_TB();

endmodule