module cpu(
	input clk,
	output addr
);



endmodule